`include "testbench.v"
`include "btn_in.v"

module btn_in_tb;
  initial begin
    `alert_empty_tb;
  end
endmodule
