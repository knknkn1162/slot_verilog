`include "testbench.v"
`include "slot.v"

module slot_tb;
  initial begin
    `alert_empty_tb
  end
endmodule
